`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    15:04:58 12/25/2016 
// Design Name: 
// Module Name:    transform 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module transform(
	input[9:0] x,
	input[8:0] y,
	output [3:0] i,
	output [3:0] j
    );
	reg [3:0] k1,k2;

	assign j=   (x>=(1-1)*48&&x<1*48)?1:
				(x>=(2-1)*48&&x<2*48)?2:
				(x>=(3-1)*48&&x<3*48)?3:
				(x>=(4-1)*48&&x<4*48)?4:
				(x>=(5-1)*48&&x<5*48)?5:
				(x>=(6-1)*48&&x<6*48)?6:
				(x>=(7-1)*48&&x<7*48)?7:
				(x>=(8-1)*48&&x<8*48)?8:
				(x>=(9-1)*48&&x<9*48)?9:
				(x>=(10-1)*48&&x<10*48)?10:
				(x>=(11-1)*48&&x<11*48)?11:
				(x>=(12-1)*48&&x<12*48)?12:0;
	
	assign i=   (y>=(1-1)*48&&y<1*48)?1:
				(y>=(2-1)*48&&y<2*48)?2:
				(y>=(3-1)*48&&y<3*48)?3:
				(y>=(4-1)*48&&y<4*48)?4:
				(y>=(5-1)*48&&y<5*48)?5:
				(y>=(6-1)*48&&y<6*48)?6:
				(y>=(7-1)*48&&y<7*48)?7:
				(y>=(8-1)*48&&y<8*48)?8:
				(y>=(9-1)*48&&y<9*48)?9:0;
endmodule
